module mips (   input           clk, reset,
                output  [31:0]  PCF,
                input   [31:0]  InstrF,
                output          MemWriteM,
                output  [31:0]  ALUOutM, WriteDataM,
                input   [31:0]  ReadDataM,
                output  [31:0]      PCW,
                output              RegWriteW,
                output  [4:0]       WriteRegW,
                output  [31:0]      ResultW);

    controller c (  InstrD[31:26], InstrD[5:0],
                    MemtoRegW, MemWriteM,
                    PCSrcD, ALUSrcE,
                    RegDstE,
                                RegWriteW,
                    JumpD,
                    ALUControlE,
                        RsD[4:0], RtD[4:0], RsE[4:0], RtE[4:0],
                        RegWriteE, RegWriteM, 
                        WriteRegE[4:0], WriteRegM[4:0], WriteRegW[4:0],
                        ForwardAD, ForwardBD, ForwardAE, ForwardBE,
                        MemtoRegE, MemtoRegM,
                        StallF, StallD,
                                BranchD,
                        FlushE,
                            ConditionD);
    
    datapath dp (   clk, reset,
                    InstrD,
                    MemtoRegW, MemWriteM,
                    PCSrcD, ALUSrcE,
                    RegDstE,
                                RegWriteW,
                    JumpD,
                    ALUControlE,
                        RsD[4:0], RtD[4:0], RsE[4:0], RtE[4:0],
                        RegWriteE, RegWriteM, 
                        WriteRegE[4:0], WriteRegM[4:0], WriteRegW[4:0],
                        ForwardAD, ForwardBD, ForwardAE, ForwardBE,
                        MemtoRegE, MemtoRegM,
                        StallF, StallD,
                        BranchD,
                        FlushE,
                            ConditionD,
                                    WriteDataM,
                                    ReadDataM,
                                    PCF,
                                        PCW,
                                        ResultW);
endmodule